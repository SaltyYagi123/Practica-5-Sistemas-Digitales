-- ROM file for the ICAI-RISC-V processor.
-- Generated from the hex file:  ROM.vhd

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
  port(
    clk: in std_logic;                         -- Synchronous ROM
    en_pc: in std_logic;                       -- Whith enable
    addr: in  std_logic_vector(31 downto 0);   -- Address bus
    data: out std_logic_vector(31 downto 0) ); -- Data out
end ROM;

architecture Behavioural of ROM is
  -- The internal address is word address, no byte address
  signal internal_addr : std_logic_vector(29 downto 0);

  -- ROM declaration
 type mem_t is array (0 to 154 ) of std_logic_vector(31 downto 0);
  signal memory : mem_t:= (
     0  => X"00100313",
     1  => X"fff00393",
     2  => X"008000ef",
     3  => X"f9c00613",
     4  => X"06400693",
     5  => X"010080e7",
     6  => X"f3800713",
     7  => X"0c800793",
     8  => X"00200313",
     9  => X"00200393",
     10  => X"00730663",
     11  => X"fff00513",
     12  => X"230000ef",
     13  => X"00100593",
     14  => X"00100313",
     15  => X"00734663",
     16  => X"ffe00513",
     17  => X"21c000ef",
     18  => X"00200593",
     19  => X"0063d663",
     20  => X"ffd00513",
     21  => X"20c000ef",
     22  => X"00300593",
     23  => X"00639663",
     24  => X"ffc00513",
     25  => X"1fc000ef",
     26  => X"00400593",
     27  => X"f9c00313",
     28  => X"0063e663",
     29  => X"ffb00513",
     30  => X"1e8000ef",
     31  => X"00500593",
     32  => X"00737663",
     33  => X"ffa00513",
     34  => X"1d8000ef",
     35  => X"00600593",
     36  => X"00200313",
     37  => X"00100e93",
     38  => X"00a32393",
     39  => X"007e8663",
     40  => X"ff900513",
     41  => X"1bc000ef",
     42  => X"00700593",
     43  => X"00000e93",
     44  => X"f9c00313",
     45  => X"00a33393",
     46  => X"007e8663",
     47  => X"ff800513",
     48  => X"1a0000ef",
     49  => X"00800593",
     50  => X"00600313",
     51  => X"00400e93",
     52  => X"00234393",
     53  => X"007e8663",
     54  => X"ff700513",
     55  => X"184000ef",
     56  => X"00900593",
     57  => X"00600e93",
     58  => X"00236393",
     59  => X"007e8663",
     60  => X"ff600513",
     61  => X"16c000ef",
     62  => X"00a00593",
     63  => X"00200e93",
     64  => X"00237393",
     65  => X"007e8663",
     66  => X"ff500513",
     67  => X"154000ef",
     68  => X"00b00593",
     69  => X"00200313",
     70  => X"00400e93",
     71  => X"00131393",
     72  => X"007e8663",
     73  => X"ff400513",
     74  => X"138000ef",
     75  => X"00c00593",
     76  => X"fff00313",
     77  => X"7ff00e93",
     78  => X"01535393",
     79  => X"007e8663",
     80  => X"ff300513",
     81  => X"11c000ef",
     82  => X"00d00593",
     83  => X"fff00e93",
     84  => X"41535393",
     85  => X"007e8663",
     86  => X"ff200513",
     87  => X"104000ef",
     88  => X"00e00593",
     89  => X"00500313",
     90  => X"00300393",
     91  => X"00200e93",
     92  => X"40730e33",
     93  => X"01ce8663",
     94  => X"ff100513",
     95  => X"0e4000ef",
     96  => X"00f00593",
     97  => X"fff00313",
     98  => X"00f00393",
     99  => X"00612223",
     100  => X"00611423",
     101  => X"00610623",
     102  => X"00412383",
     103  => X"fff00e93",
     104  => X"007e8663",
     105  => X"ff000513",
     106  => X"0b8000ef",
     107  => X"01000593",
     108  => X"00811383",
     109  => X"007e8663",
     110  => X"fef00513",
     111  => X"0a4000ef",
     112  => X"01100593",
     113  => X"00c10383",
     114  => X"fff00e93",
     115  => X"007e8663",
     116  => X"fee00513",
     117  => X"08c000ef",
     118  => X"01200593",
     119  => X"00815383",
     120  => X"7ff00e93",
     121  => X"0053d393",
     122  => X"007e8663",
     123  => X"fed00513",
     124  => X"070000ef",
     125  => X"01300593",
     126  => X"00c14383",
     127  => X"00f00e93",
     128  => X"0043d393",
     129  => X"007e8663",
     130  => X"fec00513",
     131  => X"054000ef",
     132  => X"01400593",
     133  => X"00001337",
     134  => X"f1130393",
     135  => X"0f100e93",
     136  => X"0043d393",
     137  => X"007e8663",
     138  => X"feb00513",
     139  => X"034000ef",
     140  => X"01500593",
     141  => X"00001317",
     142  => X"00000397",
     143  => X"ffc38393",
     144  => X"00001e37",
     145  => X"01c383b3",
     146  => X"00730663",
     147  => X"fea00513",
     148  => X"010000ef",
     149  => X"01600593",
     150  => X"00100493",
     151  => X"008000ef",
     152  => X"fff00413",
     others => X"00000000");
begin

  internal_addr <= addr(31 downto 2);

  mem_rom: process(clk)
  begin
    if clk'event and clk = '1' then
      if en_pc = '1' then
        data <= memory(to_integer(unsigned(internal_addr)));
      end if;
    end if;
  end process mem_rom;
end architecture Behavioural;

